library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package prince_cipher_pkg is
    type test is record
		key      : std_logic_vector(127 downto 0);
		plain    : std_logic_vector(63 downto 0);
		cipher : std_logic_vector(63 downto 0);
	end record test;
	type testArray is array (natural range <>) of test;
	constant tests : testarray := (
        (x"00000000000000000000000000000000", x"0000000000000000", x"818665AA0D02DFDA"),
		(x"00000000000000000000000000000000", x"ffffffffffffffff", x"604AE6CA03C20ADA"),
		(x"ffffffffffffffff0000000000000000", x"0000000000000000", x"9FB51935FC3DF524"),
		(x"0000000000000000ffffffffffffffff", x"0000000000000000", x"78A54CBE737BB7EF"),
		(x"0000000000000000fedcba9876543210", x"0123456789abcdef", x"AE25AD3CA8FA9CCF"),
		(x"49f14b6bf3d0e6364f86b184b3bca293", x"357947981fcd2c8b", x"0E6657D4C7FA2FE4"),
		(x"3af6de0b7eb0efa22f0210964f864fee", x"32e5ca087caf7c7d", x"F9ED3E9EB35E0B38"),
		(x"82312b3a81afa6a080d8151ba2d5a036", x"08b99f78e802b4a9", x"605ACB8772B639B2"),
		(x"7901d040d0f2710d3c5b65d19298b91d", x"5111ca9ec1fbce8b", x"7350E6C1DE34BA94"),
		(x"111e485ece3f3cd6ce5e7eea187c234a", x"225f1efdc14bf647", x"E72F58BFC2BC00DF"),
		(x"608fe310182a197d095931433def1414", x"95f9a142793a73fe", x"CD331A688BC6018E"),
		(x"67190c79c6c35b1ab779d7854a294689", x"701fc94781906d06", x"6EC55CEBC52205B4"),
		(x"2fee48b0fa96dcbd031d223b82037d24", x"eb64c15f06a40a25", x"90DE8754C132A90C"),
		(x"d5b301233199fe44f85d474a108a6fee", x"62042158c51cfeea", x"C53F0CFD97214FCA"),
		(x"f539ab1b59e68c9c21c4fb5cc12248f0", x"6c7eade673a16b32", x"9B7896223CDC59CF"),
		(x"4f0aa94c5bd4b9b5a5b2db75d6d4e49b", x"d62eb3f0d05e62d1", x"A12A1C7FEDE9C32B"),
		(x"c93320228e84c37a647e910027e88762", x"0c8608a968354994", x"9CEF3743B9E74F01"),
		(x"619454c3cd507b8be251f3ffdc679334", x"359d157069bb0711", x"CB41B9B8C58B63AF"),
		(x"266124bf1ab187a70a27f58123408227", x"310276732cedce7f", x"5C9C87477B66EDC0"),
		(x"6c47e3c425d6c879a2c67a0cc2e771bc", x"51e9c3d9aa73e233", x"39BFB6EB18C7FB79"),
		(x"94ecfaeede590b389af372a549c3a9a4", x"7b2adfbe11503278", x"3B097B1BFB3DA7F0"),
		(x"cce18430fc8e7efea550da5c605a737c", x"ca4ff15003ebc06d", x"666CCA309BC561CA"),
		(x"6afeb42ae67d75790bde22077f796929", x"1e0e41ebcc19f9b0", x"C1984BA496BC6177"),
		(x"58dd952290eaab9c529c197316a58e55", x"6559e6e06bcdef9d", x"5B9E2A3D529E2FFA"),
		(x"c9ab453c3903fd96662370e5f4663460", x"5a8808cb19670a78", x"72D5212511E02753"),
		(x"7ac956b69bff0e041460cbfd4c49da60", x"1c218ce5ef14ccba", x"1C97AFFE137AE0B8"),
		(x"f46649fad982fd9399a9143e93899638", x"feadd8df20e9f466", x"9A4A8967B2831746"),
		(x"3c674ddd02fe8843d0f0c6d1f1e6a2cc", x"e1ba30a673a4db54", x"BDC9E69BABFD1EB5"),
		(x"12f5bd1a2c3cf46422bb7ba903aada40", x"c573002cc8a1724b", x"7CA616E16394278F"),
		(x"1360e046042b0bcf1e1932a2e58db787", x"ff9a973744894149", x"C5280998044FE377"),
		(x"e8b3018e299eca253d954f56aa7a6d07", x"f45afe979fd88823", x"8990C492F1B4B8EA"),
		(x"172012211b7a590d7a8908cdd9549d0e", x"956fb84c331c35ae", x"414E46C392A26A31"),
		(x"2fb73e1bc18cf35a3b8a9b45cbfe6e29", x"24d7f62e3a1fe248", x"5F2D897491290B2E"),
		(x"2fba218e429680691f28015cb67ee067", x"8252cb89751ec74f", x"04B7F9FB38439C8F"),
		(x"5761da28ddb2506b9b088788249d2ae2", x"5f6c85c63f959804", x"DDEB9384749F96AE"),
		(x"838cb29f8d7bd80719c3a6fd5c253689", x"9737f2bdb1c1c60e", x"C77C961BC3CC5527"),
		(x"1998c53d49e178dc11a781e7c4ddab45", x"8b022c2363aff8a4", x"09B53544CCF4D59F"),
		(x"c4fb56ad583c67eb1bd13732e11d8f1f", x"1331eb75579fd2e6", x"41BC1ED10886A03C"),
		(x"c7e3f474f2d2ac33b1e29c5fedfc2d1f", x"823ce5decec48e4a", x"1EE9521A6A60F5F3"),
		(x"06d80367ba0562cdc4eca3ab4e32f69f", x"dcfdea8457833a81", x"DBFADDF8BC1D36C2"),
		(x"5fcd6b1b8f2a2c450309285b2bc179f2", x"943228311ebbe9bf", x"F31D2964D0BFF44D"),
		(x"581671c61b1de220ad41daa6ffd33a59", x"5490672f2bb0c158", x"DE5AAF2A4C8F5931"),
		(x"b2a2c3109edb3ecc676b5cfd78579b77", x"93abbc2e5b4bc473", x"92DB61DC10622A7B"),
		(x"236f3bed444c5dad5525a1b59bc99c3a", x"a1e969e6d838988c", x"D99CEA79D50AD907"),
		(x"ec8fdd04ce9bbe74642ffbf1b529409a", x"d34b1eff5f959dcc", x"C7080019A1FD5709"),
		(x"2f333f85e9c33f2e62e8f28abac02d0a", x"df160ac2ae94124f", x"F0A7716B74ACCCB8"),
		(x"b4ede70e78ff383f7732921352f6abca", x"4dc3528413114dab", x"4C76FE73ED6E97DF"),
		(x"692a6949d37b4b23aa5b8748dbeed950", x"06865629a9521557", x"F6B428D20BCFB9C8"),
		(x"85443e326facdf527037e287a78c579f", x"a96bebeed65ff155", x"06342F2DB7CE0D42"),
		(x"fc3ffb71c7c9c3af18fffc7d6c6f3641", x"57325ad60b3d0f20", x"A07AE6D3D211EDBA"),
		(x"1d34d5ed3a4e970c300e031206e31f35", x"b2b430b9f4df1f77", x"CFA061E9D0A3DF81"),
		(x"3ef63bd51917cc4ef08b9b1c72486c33", x"d1fa2b370d63dcb2", x"528BD28FDA378C05"),
		(x"b8a5f10cb60bf23abc7b51948655b7b7", x"9e959f38a1c8e6d4", x"8C024579B26E448B"),
		(x"da37c09349d389d943c3fe8f5c9a63d5", x"e4ac88f046f1f8f2", x"60E3CDC5D3832390"),
		(x"f20e2412b67ea82ec7ecfd049eb406d6", x"c274723a829dcc5a", x"734DBB62FC34B6B8"),
		(x"72421a38feb2c5bb13d32e2ffabb4f6f", x"d1c552fbe231fd12", x"F552490C8D25D5A0"),
		(x"44aa8ff29e7cf5fa2474ccb205f31152", x"41bfc541b934a1c8", x"BEB1565282C1D5CF"),
		(x"d483b24db1bf2113f7b7f92ef41b24fa", x"b69edc71ebf4ae5b", x"FF13337FC641AE66"),
		(x"31d50fea971d84b44745adcce44ead2a", x"5d11635bd2586ae0", x"EC1E67845C43B4F7"),
		(x"0a90fbada1b53857b599d353eca8adf8", x"fd62587295164e3f", x"44A42BAD0F9EE70B"),
		(x"38151e295a44c6c0b50e674d5ccd5deb", x"3626b3b25f735d9c", x"5260837012136E1F"),
		(x"32537d84ccb16f6e873ace22cb56be7c", x"c37070f423ce8961", x"7EEE46D7FE8EA453"),
		(x"0cc0b422c80bdc70615db77e85baafb7", x"0d725235641cedc4", x"818CBA3E30A0F28A"),
		(x"469979537d61e74aad52343c29f84c86", x"2bf2b707fb38856d", x"1565393029024419"),
		(x"8c4c49a2340af97381267044f49653c5", x"89a3b564c4a42d07", x"368B720F76F4BCCF"),
		(x"127ccd16e0777ed4ad8e94c134175305", x"1ece818c03f9e0ae", x"9ABA9E789072BB79"),
		(x"b70014a9369f34a692b9782b41b9033b", x"0063bb80a5dea00e", x"53FC65932191680E"),
		(x"39d3f40183bfadc32680d3727160026d", x"8db04fd9bb4f068c", x"57F77DC2B2CC05BE"),
		(x"65872d7db5117edf4aad10769cdee731", x"9441376c649ff58b", x"566137C59A72D420"),
		(x"4e6ffed4e060fc4289426c1b81478ffa", x"cd3589660266208f", x"3308D3BC08487AD1"),
		(x"16244e51d9eddd97974633934fc1ef9d", x"a3248b44c7cfa59d", x"986752795543A10A"),
		(x"a0f9bfba17ba15f917121841fcd10daf", x"cb591179181af08e", x"749F3D8769335170"),
		(x"c2bddbf219832989df7c3cde96de70e6", x"141b28f2e38b3fac", x"1F4CB195B15276C2"),
		(x"3aba99809cd39cb921b66dc72edaa309", x"e6c000c412c0e259", x"194EB845C63EF46E"),
		(x"3791ac2199cbf797c5c7a6cabd5a9afa", x"fe45292520640f60", x"07D5E3ED015BD758"),
		(x"e5887f446ef18eef01a920be388c7423", x"0f25b785db7a4bf1", x"D63C234B1D89745C"),
		(x"563201991913f78df77d2cc61066787e", x"8014f5b3716fea09", x"A4BEDB9FE8BD3F8A"),
		(x"98a83812037c74fd68193f4509713d15", x"6bb4ea06c7b56a05", x"3CE1D698086DA1C9"),
		(x"49daac7d83e006ebb5f337cc2e55f1e4", x"7ec447cc4f082466", x"9383CC9D92A69987"),
		(x"a6e033345e5edaad7db1e004ac91ebc0", x"7dd381d1bed0dee0", x"6E3A3767A4A1FB03"),
		(x"97418b7d83b8dac736fe28efae942a0f", x"75273f25ba9567a7", x"14423D2B11CC7B4C"),
		(x"7c31631a2749d63884fe65356d075a72", x"096b28be3365442f", x"1FCBDE8DA6F33DB1"),
		(x"39fcb451d7a401f313cf1cb8c21ac3e8", x"b4d1d6192de48baf", x"E5A97F334B79B62F"),
		(x"0a0acda947a618223ed38204afaa6be6", x"b7338a47c6b4c33c", x"E0B73BE8E3329E09"),
		(x"449995327b9abf644d9f11e35c7d8710", x"4e5b8335246c32a6", x"479EFAE1B0C30FA7"),
		(x"cb7841398af2aaa95832fbf4c64e84cb", x"befe579a940ae11d", x"87EF963510D1F0AC"),
		(x"2375ed803417547b908279619907955d", x"24c0b76acbf5b9cd", x"69574B006920D3F3"),
		(x"ac486bbb8d0330ea96de0c3d2dccc3ad", x"54896e9209e73daf", x"00A76968AE5EEBC4"),
		(x"b6484d7cd0888593305e0535e37d8105", x"f96604b9488fdbb0", x"A44EF4A4065E4FE4"),
		(x"b93e71fd773f890c788f7d6276793a5f", x"d863c5c0eb0326bf", x"2FB2B566CC4E4A01"),
		(x"0e8a74f9e9470580d94c86cbf2e5459a", x"75deb76ebc60189f", x"9E4EFFA4C73321B6"),
		(x"80527b4508993be65d6d439226ef86f6", x"2300ccc18615ecdb", x"4D86E635318778D4"),
		(x"fa5bf1026a7fefd10a3a5f8614a20204", x"d08716a5149605e8", x"149AED96296B6293"),
		(x"23bef41171005d769346e6dac4bc61cd", x"7916ae8da206510a", x"EC6172BC566DF5BB"),
		(x"a6da3b97cd1f77310441941b8242d777", x"bb68bf66faa6bca6", x"B573EE3B6AD6015B"),
		(x"8f481ec4f1ae4a4b9be004336654b73a", x"57361510f95d1036", x"02406B396804663E"),
		(x"e83b235aaa659333f36f55eee0ef476c", x"92be219174a1dd3b", x"A13F4002CE86F70E"),
		(x"2d9779a1428d76d5a987344965b6f088", x"f78f4f2c57151b34", x"8C509C4980D06E22"),
		(x"066fd0d31f667836860cae04982c16a1", x"a35c27c6bf34b52e", x"E1DEE488BCA84289"),
		(x"99adbca480e7f49aa69cddbe4c8fa8f8", x"e1b791dd84925d5c", x"BC4798CD5D4653AD"),
		(x"bab3c3525cbe288dc319bb8593bac290", x"b1454dcd48cc0892", x"33BCD18143B05A02"),
		(x"05bf2eac7341fff28885363e4dbaf4cc", x"4176cc193df9c494", x"A0D4C12F782357D6"),
		(x"30d448c1da113b7837b2eeeecd7d5a94", x"8ae6424099582273", x"CDA3379A073C35E5"),
		(x"fe55489598b0c8bfc896840c275bd0a9", x"6940836d02172da8", x"C68C0FE0D92AD1BF"),
		(x"90fecfa28d6e7ba1c57c205a92003ef4", x"56be4022548aef70", x"223FDE155C4B4D22"),
		(x"cd8ff07d15815a357b0d51f468691117", x"23d7811bc514562b", x"6779A36928096694"),
		(x"6b02d714629770d358d723a2fd8c372a", x"ba25a3de04a25918", x"C0341FEB94FE3012"),
		(x"ad90d6d7d5269a1b08e413e7b5e6c443", x"293e3d712a6f3464", x"A35954FCE2B33B5C"),
		(x"510a9cd3c345a03885fb507e5dd6f7bc", x"24068e9139d4f509", x"2CA8C175AE084597"),
		(x"446e21d8c5fc5675b33ccddaabd11b22", x"aec6cc12783534fa", x"899F32556056FF18"),
		(x"76a0a0e1c64779db055926411dda3148", x"65e3286d2f59790b", x"1054C47949FA2348"),
		(x"bb1e4c3f62dd7cf5b9d17130450d131d", x"9c6b97e971c17f26", x"667AE666566FBDE7"),
		(x"4afba7648198636aed1c744e70a6b1d4", x"3e5ad72acc0e39a6", x"13D4CEF720174CC2"),
		(x"4782da1885263e62a61fe3b3c42433da", x"81c87648f0e91dfc", x"0735BC857691FC58"),
		(x"cd05048cd1ad5ba8ed31b4c514ccab97", x"37a555096652a7c0", x"FC3AE60619D46109"),
		(x"883c5bba6d20ce221de3397389eadabe", x"92c1b0bde6b01305", x"99DFE2174B88EF81"),
		(x"14967dfced514c0163ce47e8ce019e3e", x"0cb764280c96bad6", x"6704A082536A9A15"),
		(x"546b669c4c24bcb52474342698ff4458", x"ba8625d7e62b69a0", x"A5E52908A5C06811"),
		(x"c374eae292aafbc2deb0ee9f79e2a248", x"a2d33bef4b81aafa", x"F48E7620762B65DB"),
		(x"c5289f515278571110247901341c5ed1", x"aaa40fabdd7430d0", x"AE2DFD6B4C1E0203"),
		(x"bb4fbc2b623666012490910e2fcc3948", x"de03dd2d0ff134a7", x"19001847EE53460E"),
		(x"93538e6fd17b4dfaa24fdbc383fac8a7", x"64a39a2672ac8301", x"5BE249DDC7BCD9C5"),
		(x"7f496ccb8392ab7536a19134ec31455e", x"5da90b935ee081b4", x"F610CB2AA44B5B93"),
		(x"e68883ee29b45a8e52e7be7c926e15d3", x"84821f6672acc868", x"87F5B0484B269B0E"),
		(x"d8cedda03977d8925f4bd18023a54244", x"303a138e90618bf5", x"3072B00DD75FC6E8"),
		(x"cb5bce9e8761e21a19f57f9ea34abe8c", x"50ac0701cc70e1d1", x"8A0FFFA8D5CF0A9B"),
		(x"cbfe2b1b75b77de3279181fd44fec543", x"3b93f810a770032b", x"1185276CF6EA9149"),
		(x"a45cb587fc6613805dc4137c6c2cba71", x"a7c4c7aede5b1a53", x"4D91DE0A32E6A775"),
		(x"aca3e346dcd090aa177b1145e410953e", x"8fa9164ca5a6145b", x"B66D3CF1104C340C"),
		(x"07b13f8512acce90391360cac3824ffc", x"05cd8c97d597f6e5", x"BE52849D23BE4E1C"),
		(x"5e973ba9d39aa84dee84529eb686180d", x"1717cb80a49c127c", x"DE40A8578675A2BF"),
		(x"ea26d7e9df0862264d70ea93d192b77e", x"81574dc2492e02b5", x"82F105F0C210E223"),
		(x"e115cb2d575fcccbf94f1f554e27a5e3", x"cebd0503c6426077", x"F57D5BCFC65AAFE9"),
		(x"598c143f2f4cc43daf7c3f37e8ef04ef", x"aa9295ba49739a2f", x"81023116F86D9F44"),
		(x"99dee23ba3e008c226447b109d00cb98", x"061d0a3f7df7d42a", x"25A9889F5ACFA296"),
		(x"e921c5e72714e61f0f20eab99d7eb86f", x"33461f09ad0dc7d4", x"1F8005EB8EBFB58E"),
		(x"01df59483658e713ee0d862e79078252", x"8c35852226a7c707", x"F41ACE1DA57D74D2"),
		(x"95dd63aeca78cf5589b74bbeb81f38f6", x"70b963e6b45fade7", x"3613F3D0F1BCA470"),
		(x"93b193ae701db1077513153137bd3ee3", x"aaecf0b6e5b1e974", x"A662D2908275D92D"),
		(x"f390887e5d4e2ec4a8e6bac8845dfdfd", x"62a78b2827c73465", x"7C435B3E5F17B233"),
		(x"c730f6bed1af3a9cbf319d253a80298c", x"2ab86981ddb196f9", x"C533C9CC927F35CC"),
		(x"3783abcb194f9f62aa022f0b43ce5d51", x"f93efa43dc3ff33a", x"76E7A764F9C73718"),
		(x"146b468d96ffe542b988cee15a6db034", x"56a150f2556832df", x"0A19AF10DD3FC8DF"),
		(x"a31d91ebc493791bb48fe0c94f7d5aa6", x"68fb5d416a7908a8", x"48C47135B830E862"),
		(x"bb6a57db41264df52def9a5ed5631170", x"7b79c9216078fb96", x"1C8C95055A6C40A1"),
		(x"21e9360db3420bbf55c6c339e187b847", x"e82755e0c688bd42", x"0CF3EB1C52864425"),
		(x"10a66077a9444cc2d9f634a20b052c99", x"3a28d37e4374a8f1", x"922D330B9004FD77"),
		(x"23a06f1daca762086aaa5cb1d2931b44", x"5fa33827338eda63", x"27200E537F3DC3DC"),
		(x"7fc73c1e4bf8145cfada9b1ff63f517f", x"b5a573bcc02d2fcf", x"BA125A6108D474DC"),
		(x"2d6d910f8f0b43128c59766db8868b9c", x"75235bb776dd3c86", x"2072BC24E906B1D4"),
		(x"03929f9ac21a1eef7cfdfbceea4baae6", x"b8e9beb1ada32e07", x"919186D8080BD063"),
		(x"2703f9bb07f0c94afaedcbd86bff21b9", x"9603da31ba67ba41", x"2491E02F2E450161"),
		(x"89685933a008de16276ecd6ba5dc5f81", x"e7ded24e6d875747", x"F49F87F70607C77E"),
		(x"c53e3ce3df41da17a7b25d7d490e0303", x"de32c498f658c894", x"6E99747721C76EEC"),
		(x"ece64ad2585d3497d2732b14a2e0fb3e", x"4b63a1ca25fd477f", x"8C6C6D548D8BDC5C"),
		(x"baf8a62719f428df9cf714af08aac1cb", x"f263f385998227e7", x"B073B9D30C708CF4"),
		(x"d38acb6e95f0c9d3f5b0e7f4dce06031", x"4e577d643a49293b", x"854B313670A52821"),
		(x"807df259219a029f69f17f4d4379a6fa", x"4bf68830ebe17fac", x"7019EAB5832F7C0C"),
		(x"106f6716f9144e22320a51fd8b1c54f2", x"26218a5385d95ad1", x"5E10ABADFBAF1A90"),
		(x"6e93fe45337a69233eafa7fc7b75df05", x"2aa8648941918e42", x"6644A338D9012092"),
		(x"56c387432ec966b4751138a61e6a58d8", x"84cc347d407509a4", x"C632CBB29F3473C2"),
		(x"5312b796feafb98f4002e2dd9519a06c", x"76ac1631b4cbaecd", x"C9077F3BC5F18124"),
		(x"100e113fc756d5978a8bed79cce09f1c", x"723ef33c9426f1a3", x"7A3FCC17909922AF"),
		(x"662b823a62b56675aa9b6b6d55d0b85e", x"502a4b1178f90ed2", x"3D08EDF18FA80962"),
		(x"e82bbeaac4ff8d6aa035d7bf34a6be0a", x"6236c831e685fd4d", x"711C01579F4E111C"),
		(x"1fe0c657267f7ead05eee0f27e5f1b90", x"718d14c4216c082c", x"E50CDB1453C23375"),
		(x"0fbea26154dfc7701d4f139bd309a474", x"9fc6ad5d22f0fe7e", x"1BD5CAEA5339415D"),
		(x"6bbdcdc9ae11094bb7fb22524c4d2fef", x"b1df2024c18bbd5d", x"E5769DB8BC8F83FC"),
		(x"fe93288fcf1a2eb5fe2a3daac8e5b2c1", x"cd1b50314fbe69af", x"05CD57F649879CF1"),
		(x"6b718765db29f577744769662df238f3", x"e85cc7f880ce3251", x"FB5AABDBD8664788"),
		(x"f09ed05810707b422cc28b17ff16201b", x"39647b243e0f2d41", x"85C3AE0D3463DE5A"),
		(x"65ad8eed5770dbd2918d2de25b1fc2ee", x"b065862b36ab5681", x"6830594DD2DC178F"),
		(x"075da0aba24f154d098366e9ea316230", x"0f5419c585f4c483", x"AE9921B6441FB069"),
		(x"9a0e2dde0b0823039e82714014d810e0", x"5d56e5e8853688f9", x"E57F20B5848FDD30"),
		(x"3bd9b6dc9dfd9adbdecc5e18ca4a8540", x"f21edd3d96566848", x"AF481A5A2CFE1B68"),
		(x"04122ed9783eb51fe9916f664066fb0e", x"d392b8b6219b7b37", x"2C4D842DC1E11216"),
		(x"613be1d2180212001e6839ec02df7228", x"313c2106eb35bd93", x"EDE0C066C768953F"),
		(x"d05c186e6f3570955fc02a31ab17de52", x"f0ce0fedf85c30c2", x"D3CF25D4C1D747A4"),
		(x"568c135d0779fde16b73b2ec8797e62d", x"dc59d9278ad1991b", x"B1A3D63D2EEEACAC"),
		(x"d9888dbd2b9d007c93fdcb83f1354f78", x"c2e6df07bb8f3f6c", x"5C2BB0CC1BCA170C"),
		(x"d6192a700ee126d8bd5dd38b3f82c1fa", x"3d1418f6caa9a42b", x"761EFF64D1AF40FA"),
		(x"a17b0e5b20756c609b8a5a17a29c5e26", x"05fe8898bf6a7828", x"588A39CB3B37ECB2"),
		(x"9531bb47dd1cb9f73dec2a718d30842a", x"a24680fd0dd49eae", x"5923F5726CBC3A85"),
		(x"bee3b41ffcf6efd635c16b380673c73c", x"3649208c2f5f4187", x"9B8730DDB29FE046"),
		(x"dbc0ed8a7e498a91bde532c9ca4ea805", x"79ca92564684672e", x"046CB62DB19E2E9F"),
		(x"a18717b54d2a629a6adfd553cf5385c2", x"09420ade4eedd2b9", x"B427B1B793E64023"),
		(x"c86d231fbd2933bb8d8a73c22582205f", x"1ac25a406d68933d", x"342161F50E96A718"),
		(x"a7d81643a9f5d171c927f4cee57a0a2c", x"bc9eba2db74b8631", x"73E42850CDF890EA"),
		(x"8aec23553c65be70a03801cce38eb50a", x"a1dc23ea46a37c96", x"FCED870A93B4E3D9"),
		(x"a1c9ce587ae86d1ed61349824f6734c1", x"d00eae97f8661d37", x"8505E6758D0D7FF1"),
		(x"92f9406eccaeb602737192c607792403", x"4d098b000945118e", x"43178D6DC74014A8"),
		(x"77242c5caa98be0af0567b0ba8d5c8d0", x"755df56806ce14d7", x"CE3D1D51F8111CBE"),
		(x"784e64771041babf397d810f5330037a", x"a381f9a68536731f", x"30F35A54045EC738"),
		(x"ed7fe425288293b16996c2a6217df0b4", x"8379760a87e6905e", x"1071C05355918A5F"),
		(x"ef50c820624357b553a0fd50c6308a93", x"39a017f54d668a3f", x"D3D27F72CA0A27E3"),
		(x"6c7d77937710599a42954b32785ed533", x"2dbce8012996b8ac", x"85EA7F5DCA3D4F46"),
		(x"8524ea8a6b3123c7052c6e7169eebe9f", x"0a6f6b6a18db97b6", x"8ABB61757AFEC706"),
		(x"417160148fa926983c0e5ead0c839369", x"60c20c43580915ea", x"8DF81774464B2DCB"),
		(x"f9acfdff737288b24af697033e7dc87e", x"79818875caddca4a", x"A36FA11F5831A202"),
		(x"08ed04eae86124eb7b003eb663f4d4e1", x"52b064ce4f10e4a1", x"21FABD7CE7CDC609"),
		(x"308ba4f99260d4b892b2ecc42a1f19b3", x"8d987bddd5ae2310", x"0C65ED91E0884F6D"),
		(x"12f38d3d77aead3763a5b47ca033f453", x"3bcb9ba261f1da29", x"F334A71E4AB3B1EF"),
		(x"cc693b2abf09f52950bfa4a9a3113577", x"f0aa8f6bb1f52c19", x"AC3E5B32C7E4BE96"),
		(x"2107515d55016928b77fe7c17922e37e", x"d207084de6d00ac4", x"A172D86DBA64723B"),
		(x"a2bfe624f2e48f49dc9ad8be42e0e16c", x"b2779b97ed22dbd8", x"F5A7DF8DA0EFD8F7"),
		(x"3baeaad06912a20e0c2078f1a969216b", x"b8eb9313a8bef417", x"5B6BB5D4166E3E9E"),
		(x"cf04332082deb3c5f115cb85c806a5f9", x"15e31a9f43ab6514", x"C3B0CD5B9BACC8DD"),
		(x"9fd9f65164507848a1e183ab21de1bfc", x"028c4c8331fcccd4", x"1BC16BE518F4B110"),
		(x"cbd09a8926d6d40227957a4540f3b941", x"1cd128e262ca1518", x"A6FAA444C44CF0A6"),
		(x"c52764ac5004e214155b530dfac9b493", x"e50c0937c7765119", x"12E1EF47D2FA4AD7"),
		(x"fab1079d5f95ffad95c222ff47f91607", x"3cb1a500d6a0f0e2", x"6706DC8DB7D02CA9"),
		(x"35429dfadb35e4292acd31d3e1007c2b", x"06729d64121eb964", x"489D9CB66DA32CEF"),
		(x"f897ceae978046374439565c36c6665a", x"10d49f92aebb7a04", x"1C2226950A8329BE"),
		(x"19da1dbd5a2f7c6d464b146e2e17ff91", x"83704565fe99d80a", x"B6A43BFCE4DA81C4"),
		(x"456b6e0ec5cccfc478011816973b8491", x"0b7369e605ff167f", x"0C5C4B748A46F58D"),
		(x"844bb2b28694a0d284bd9e68ffa3b0c6", x"459dbd23b0107d6f", x"B65A46C6C31EE6A2"),
		(x"0a901c0c40c2a1dc7c6a1b202f0ced2a", x"fc285ac86f84e5f9", x"542C0C47BA052B2E"),
		(x"fdd1884e44df7d4f42b9e44df1b6b9d5", x"4f0e4fd16aaedec3", x"1F8F1DBA93218DC0"),
		(x"dc5a1154c4be341a7b0d7aa5140c2676", x"de59d944368d396b", x"FACA72AE61E6BE1E"),
		(x"a24df223e3b2c3ec89a1694c69efb72c", x"efc7de9c06e4b54b", x"9E88FCF35ED7121E"),
		(x"e819500c96aad7638645f6d202ea75d2", x"0a38a7ffd1e6c995", x"E44D55FD4DC39219"),
		(x"34d6676c93cb2829e5e45425d465930b", x"c2fcf5d0f37e3bec", x"3AEA8E1E90357A29"),
		(x"80c24139ad49b822bd596fecfb2440d0", x"e860dc21547395de", x"5B6D8867F121285D"),
		(x"4b210300e6aed26874738ee65dd18a20", x"920d13418356f1ab", x"BF2B7BA6841E730E"),
		(x"9ec1836e963effb8e5e2a3780759e9b2", x"1eb21050e7302a6e", x"ABD1CD17F1B166A9"),
		(x"83251f8536359d80e7366a03171ec407", x"cdd17e397b88b114", x"D9B8C4633FAE799D"),
		(x"3a49f8014b8e61e4aa090301e604b54b", x"17efe2cd61673404", x"D02DD8B29B153735"),
		(x"bc7a30c9ad9e14b084a3a3c079b427c8", x"e44f72f2fbf7f937", x"7527FA22952976E2"),
		(x"2e56351103964cf5d1cafba7e02ba4be", x"2d435bf179a799f2", x"D6555C16EC69F47B"),
		(x"059bacc6b77c1088d97c04c8157d3f95", x"965115f084fecf55", x"FC2CFAB49A624558"),
		(x"f336bb0b9d27adc1810fe8d910c00ae5", x"2def53e105f3d7fe", x"49BDBFAECB8ADE06"),
		(x"9f2d29f9539a73d93a7625f903364fe1", x"82c746fb740a4219", x"5DA1E6E8F2902572"),
		(x"4b516904c12d2cd00d07ab3394cc6b2e", x"a0510693b9dcb2fe", x"20CE912D2CE1B099"),
		(x"976a6e3b88a5936690c36193b9afbd81", x"eb83d8543337c3bd", x"B16F4D053DEDA9FF"),
		(x"197439b2be2065bd0173f4caad8b7c09", x"d6d0890d65b0e365", x"DA8B0A00CB3D6333"),
		(x"5a9d453cbd5f796deac78bee3b20db89", x"4e58f62a4f57c4a1", x"7736F07F87C3FCD4"),
		(x"f6f615fe7dba7ca637fccead6d8a3a75", x"179149bd3038d5b2", x"8E8C5A440CE4F17F"),
		(x"7526042e580d1f19f40416049e377762", x"539599014289e12a", x"7E24C2FEA80F83EB"),
		(x"a9e1f5f8e0ac1ade3f39159890366e2c", x"c40eaa2efe6d1fd5", x"7092D26EABDFE01F"),
		(x"cee59c613fb71f8a065042fc78ec0b3f", x"558a09ed001ee8b9", x"D782496E055EB798"),
		(x"80cb4b44d29184089a6c52c7426812e1", x"a04cec254bbe5819", x"FBA59904C8A5228F"),
		(x"4dd7e1f2fb7dbb0c7ea65e9b72437e41", x"aa204fc752965388", x"25A25977BC34F821"),
		(x"68d01698545d674fe316536c2a6930c5", x"e07c599b223a44ff", x"A5F09373B06FBD08"),
		(x"66395d8161809121ecb944bdce19d9ae", x"0250abb907d7a82a", x"9A94322B9C11D10D"),
		(x"d4aa85bea88e2b52b1439859e6d7bef0", x"aeecea462f98c768", x"3D4289080B0EF625"),
		(x"e3c85da200604560dad396c3bbecf625", x"040d13cd01c93857", x"4AAF43FBEF374F73"),
		(x"9d9794cfb152d6bf553ae6faeec3929d", x"d1981b33257b1b28", x"1D394F9EDB825C67"),
		(x"03f8e7d71e5556043a0d2a3b3666e0c3", x"8bb963ad46937904", x"E952EB528EAF0672"),
		(x"603afc19a0af905d3b230a4b4244cc46", x"c5584a6ef08040aa", x"714783A79E7834E8"),
		(x"751aaf23db15dc864e3af009a63b005b", x"5b8b43f16c386fd3", x"6F6AFDF1D72358E3"),
		(x"fde1b1bc256ec67b17acdb42e911bbee", x"f83eb3893dfe01c8", x"2BBF94B4EA86A231"),
		(x"4cb77c13dc8bbd05df147d0421389655", x"d0783b4bbe6a9cc1", x"67D2311BC8231AD1"),
		(x"5ab56565b0f64a4d95808766f7d39d47", x"da1e0287b95c4944", x"D63EF9FC15401616"),
		(x"1a1ff485f9715e8c67cbd0c6807b1774", x"ca18137ad220dfe9", x"AE51CB53077DC610"),
		(x"6e03acc4871fe4258d87bb47802b1a1b", x"40b1ae9377893e37", x"B46C00CCD899BC1E"),
		(x"6f9f6731d359a65d73d50a0b82a3c8ec", x"4f012b0e630874ad", x"5DC8A322E270B20A"),
		(x"040c8276b092608aa6b77a1d324b8193", x"2f83f49a59f42404", x"CBBD5817E81F752D"),
		(x"bd2df955e2f028078bc4aacbcd613f21", x"812c4ce07661d037", x"F46522454ACAE535"),
		(x"5743f5ca45c053ba6abcedffe19fa46f", x"332f2e66d9cc2b4b", x"DEC3374940A6CEAD"),
		(x"d1f60cfce9467d711b1e5fc816a9070c", x"fb4e3ef0410a5cff", x"035760F0F99BAEB5"),
		(x"7fe669d9fd567e1489e6ece5b92da09f", x"89b0620140de2547", x"2CE04B6D0BC119D7"),
		(x"04372797a598362eaa3030290af4bb14", x"2f463acf3e6bdfb5", x"29DD4A3189C678FC"),
		(x"a1a2230e992b3c47ed951d8732d21483", x"fb4c6c19285c9836", x"FA6622FF8F752B16"),
		(x"f6f2179ac603a59226b9742a3f84f768", x"89ec383379901012", x"D57549ED2E22F29F"),
		(x"2ab0764f3c7b32f0ef2633041936c155", x"982a58bdb3d487f3", x"CB77DC571647F453"),
		(x"92a2e686fad3422dc0892cc61dbc5bb9", x"1e829fdd6a6e44a6", x"C965BE21C16B994C"),
		(x"df2cd5fda92d67146ff33b5df06611bb", x"ef2103f6b216668f", x"A02F74793CA614F7"),
		(x"9cfc3d0d22c231bf863c167b21fa14ee", x"9ff94fa934cde0c9", x"DC702CD3FC356E49"),
		(x"ac17145ad0ea12a0d7317f3610d8cd41", x"f81e3024a6386f1b", x"508FCBFF4D427329"),
		(x"4fe57c25618b1111765ffce718a95f22", x"dea94c77b1412002", x"558EC587465A561A"),
		(x"95c393a895e738cf24360c397bee011f", x"b7047c52b3d94069", x"D0296F7113A9F5A9"),
		(x"c3184ebbda9253ca0adef6205998a3f5", x"95f8a4a790ef7f18", x"60FBDF34A9AC5C81"),
		(x"80a7ae99f48fa8b20a9e7aa849669d7b", x"8054f751407ab6ab", x"19DA6C7FA9099943"),
		(x"8383418ad6a6696a045e5cf4b891614b", x"d0f2423ef14e92e2", x"497495E9907EFC8A"),
		(x"48fe37cd9cad56396a93284cc9d9491b", x"7b4a07a8b501b560", x"9883D667572C1200"),
		(x"4510a7638b3c0c822a573ee75d66abe6", x"bd295b74b0894e62", x"2A2B00631D4290BA"),
		(x"8dc5757ef44ebd1c521faac98e918d76", x"dc4d418f0d10fb8a", x"1D2DE9085EAF002D"),
		(x"4a5d6f189cca70894178b8f1a4923022", x"b2cb93af713cb80f", x"AB5114383672FA9E"),
		(x"4874261fa6606ba03c16671a2a3a8a99", x"aff5a10ab4f87dd3", x"F85D10B04CF31C6B"),
		(x"eb0c42d8c62a5f8186408c65ad2efb4b", x"1fb967114ca12948", x"02C9640A9DA45EDA"),
		(x"d19c1eaaab11a5f830937a55621f8317", x"db947d5bddf6825f", x"F9B87B42CDEE22A3"),
		(x"0ebeecd567aedc91a1d80862eec66616", x"b30652acfcb3a42e", x"52D4EA91DF4A30F1"),
		(x"7deba9fa55d865a07ff22b75e6777fc4", x"9e652099743c2da8", x"923C4F3DA13C4BB2"),
		(x"6cd9cda5450ec1fa4662121d298c5899", x"0e096118c121a3f7", x"EF66EF37C9E67E04"),
		(x"79eb57c4e59c7e9e83a27482ce28d747", x"9b13bec9ac7661d1", x"F05C482ADCDF255D"),
		(x"aab84dd94e3431e5d66cf1bbd25ec4b4", x"d98da6a7dfccfaf8", x"BEEFD1A98590DAA6"),
		(x"7070637b20cee906ebc5db1e883b20d4", x"500021978043bb97", x"83C96E6FAAC74F99"),
		(x"675779b178873c0caa099602c5c96996", x"e249ee1e9549f054", x"1CA85003A1620C0D"),
		(x"10c51d516faf99d07c1185929b02a425", x"165f19a2072639f2", x"57F9A0EE810C6336"),
		(x"a91188c4d75d123b1244fef529cf84c8", x"592013625ac55327", x"5C60FAFAEC97A492"),
		(x"5a6a57b1cef0ddfa889a15e07b474f04", x"1744f1eb470c5bfd", x"B25DB79CEF65B088"),
		(x"9a2faf0d628ce022fdb80e7afbd05003", x"26e40aecde753599", x"007CB9D27D1DDD8E"),
		(x"f12da3dc7a39a397b6f470981d745cd4", x"663485844452b3f3", x"DD5BBEF92BE30404"),
		(x"76d40e6702d2425f53be19d8f1bc2f77", x"bb701fe2784122e1", x"FCFDDF7EC09D4698"),
		(x"faaf0b93d47565105210a99776db338f", x"6db08471ba012bc6", x"8389B6DBA5AB29AB"),
		(x"f91c5e198b919211382c710a57e5ff82", x"7c035ad3c5151137", x"0FDC93B431879237"),
		(x"963c265efed3ad380c2ca2cb0a9370ff", x"facfe9fe611f42c4", x"5F4BFB45003AB423"),
		(x"db334a02c6669f6899f352c2d29515d8", x"7818946225eea7c5", x"86BF8B9E76723E0B"),
		(x"8f18a2030ced5cce75f11df56dd00d9d", x"a60ad860730b599b", x"254D5A6AB771C36D"),
		(x"4fb1bd18954fecc655455978331674bf", x"3ce1911908151c32", x"A6458A99E9DC6253"),
		(x"ef1196ab5c6721e4cd1c6bad4bb89c88", x"605d8028ce17f932", x"84885C21E03083B0"),
		(x"c699db175cae70bdb082979fd2caac72", x"4cd6846d71af5931", x"6B61155912A7812E"),
		(x"43b391438f44619eee2e5a2fa1e0c30c", x"9e02b4cf8c5413b7", x"A7D7A69A8DD89BDE"),
		(x"77d23f59fb19cc4245e5dc46c891c840", x"8385bed6a287672e", x"2546C6046ECB8800"),
		(x"73aa5800650d12a7cd065aa8ce7c4564", x"e316c98dbc3d5586", x"A619578B53E68973"),
		(x"768c47a698d9f8b9dfadf70048d9abf4", x"923d8bbd718298af", x"133D96558C0DFD41"),
		(x"bd1e9bd96b2dca1cca513a4b5de2c336", x"d80d9272e57003eb", x"7B40B912AC490F0B"),
		(x"6dc0e542c68dd98eb6e8f6d405da6599", x"bd51f3a1cd4c027d", x"03C498F37C7F8D65"),
		(x"59306555327920b1f3dff2f8f5257b26", x"59df7e324837ff49", x"9CCE751EB42764F9"),
		(x"09da31b76d0be99fbc19977bed9552ab", x"93a7cb439122b1d3", x"D67713543F11324E"),
		(x"616ae162e4d355f8f8648fb2e0bbe2b2", x"54a1c1c9cb329762", x"B23F21AEA463F3AF"),
		(x"1c273d6a3a28bcf1ebd63b437f6af64e", x"a992f8f5ea165e7b", x"6E7A503B0FDF16F3"),
		(x"a7fd40ef60b3bd035a85e1330eb5b37f", x"d53b0b1030707a6e", x"C17B3B8FBAC49F81"),
		(x"aaaad78e180096067bbcf84acda6a818", x"24336cd587901a28", x"A685B6002D540A22"),
		(x"604150f9c2d19c654cde1168d94ab073", x"c5f9ccef7b6f546b", x"0FA26B66E9AF8937"),
		(x"2a5dafd1d21abe4638b1051a5d61e928", x"252525491aa21e82", x"F0A24355F815E897"),
		(x"e8b8bb33a15ed46b8050ed16d4303c5a", x"cc938fc5e55810fc", x"BEBFE1032E548B65"),
		(x"6dcb663ca54f23dbe6114649f63bb89b", x"7e1861ed2c5b9264", x"2B1172E76F035658"),
		(x"591b5b2cdf3172e7cb3e53db1d4a51ff", x"a4cc30f04a7a0a7b", x"09C6CBCDAF54A647"),
		(x"80cb2a3c12cd503ac354c391adad6a46", x"b54a028ce8c0ae1b", x"E6B8C726ED6CF20A"),
		(x"93d7015d7e4721c392834964fabdf75b", x"c0eda37973766186", x"4E138C709CB31F7A"),
		(x"d130a72eac9f8ab552bdc6ea01e97887", x"d658c09fa6921e61", x"44CCEC9B65294A04"),
		(x"972a92203bbe98c2ebc92177b1b4aabd", x"03d79be1fbc9bf5d", x"47684CBDB263037D"),
		(x"11a26f20c37d7cf023454939b020166c", x"78f56b06da33dc6a", x"7A97B495D53EE832"),
		(x"b22e92a8e7fcf73b85a4bbbc016f4137", x"966a0d26dbe7391f", x"89E1E982E5B69E90"),
		(x"436de05706af55098224295c2928b411", x"d86ff4378ca43f81", x"3B3BCA824992D120"),
		(x"6df546c4beb9620fef33a5bf7c3bdd29", x"ccbb4e4dc26a4d64", x"8238B165FA6AC4FC"),
		(x"86a5656d236a33fe3a12784ccef506e0", x"e4f6737fb01c441e", x"981FDB9042147C5A"),
		(x"b3a8ced4a68681c1e30e477f437a2d28", x"bbb26534e7031796", x"13DC435E8738C296"),
		(x"5dfacc7043c065559a2704100654df9a", x"93c91328b8f78d93", x"08908F7418CBDC4A"),
		(x"64cdf0a08af33cb0b219267b33b01767", x"9dc15ba509920340", x"5D246ED698043FE2"),
		(x"931b910f182ed40abd38764db601c30d", x"0d19a672c4d706fc", x"440017692754C271"),
		(x"28f36e530004fe95b6443852a7e0b8af", x"886f9c5a0efbf28f", x"190409CC8C0ED4A2"),
		(x"abf0a3c818ae160acd1abe133b2da625", x"420ef9022337f4de", x"EAF3E37C9AF8415C"),
		(x"badfccb4468ee01070f2d79e20816ebe", x"249a54335e799d6d", x"507FA9635DB76195"),
		(x"2ce172521b02c1ad1e0ea962c0de8f04", x"4dc575af18fb96d3", x"63D5CD57EBB12ECE"),
		(x"d929ac51ab6fd9a40d9ee1c0b54f9fc0", x"da3123b261106b88", x"1083C73A0B02D251"),
		(x"6b78c251a6247816e9421b01a115f25d", x"97d16a454f69817c", x"7EBB647596173D2C"),
		(x"a813828cdb4946825a61b7b011f0dfa7", x"2b2843094e72b992", x"763277B6F6DC9C0D"),
		(x"65f58a75acb1a83c3f6cd19756f24afa", x"09c11801aa5d8f55", x"C7CD4C4FDE1E7D24"),
		(x"65f767fe5ef924bff8938a23cdcfddbc", x"01d997517870293e", x"1F5A508D2474272A"),
		(x"f26d2f671556e96a4a7a7dc38198df2b", x"69b2e28e5a366cd6", x"F0B1DAAADC2C1F64"),
		(x"ee7ea2c49b1161106e5d2ef6f76ba38b", x"39e8332e2bb0de42", x"01A480E5C20331C4"),
		(x"aac299d7a62867f894a729e7cefdb5e5", x"65dd6ed64ea7270e", x"8AA784B929228397"),
		(x"4c1106a7a2b93a313fb610c7c1831b09", x"d2714529a0f93980", x"DF41EA046C1434E9"),
		(x"5f466f326218216ea09e07bf4b8a051f", x"6cd6efb72c2e8648", x"3A9E677BED29FD5A"),
		(x"05a52db1fdaff4d0be8ac393443257b3", x"df2a975b6568afd5", x"9AC61622659BFA7B"),
		(x"00c7bb5a95fbc9a8f9552e54795a5048", x"96bdf54f374e3c9b", x"F3D68BDD3592A6FE"),
		(x"cc18e7b6351f12aac482646d6970dae1", x"46f941e0684cb010", x"45C5441091BCE078"),
		(x"dcca8518f3b1d2bfb8182e86c69833a2", x"a4e42f17d715022b", x"86B9DB48E1A867D7"),
		(x"416d27ac62881dc9bfa77054a949f378", x"ca1b34faf00a0d5a", x"A382F8D48B1CBC87"),
		(x"be23f6d25b304b98798fdd47baa55249", x"916d732bafed3cc9", x"22C898C44A6F6137"),
		(x"78cb4dc4a280bb61b1471456241d740f", x"c1837507a823d37f", x"B57B6B58EC66BFF0"),
		(x"a09a7ea5d014c5e972c77832706caf77", x"37e52a261cb45567", x"F1F528A3B2BA9B5B"),
		(x"07d7d47b64935154bee7e7c8f3f4cb9e", x"4c177405185d7577", x"7FEFEBC330212663"),
		(x"ad2ee4f7ea810ceff15dec8790c0b988", x"c3c235f66146b1ba", x"EBF6F5261595BDD9"),
		(x"979890fa4c01a14203f7ecc4d0981d89", x"53b2bd29ca8cd517", x"FD82327B263DCAD7"),
		(x"e11db3f8cba464faa3277fc1ec8c1501", x"fa57e34f89fc1e1f", x"89F3E70808C7F17A"),
		(x"776537cb473b06d443899b4b2156e6c0", x"28c4e8b21117509e", x"E6A357747BFFE45C"),
		(x"594579d3eed3887abbfdd965574fc56f", x"6680aba3cac9d0f2", x"060ABE03C73583B2"),
		(x"0e0a8eae20c1ca4c8edd4e1fab5895b4", x"0df9236fdcbfe26a", x"90A23F9210B2CD1E"),
		(x"c11c86e83de1633d684b3dd35a36220c", x"48041e797a278a27", x"BCC8920334DC93A8"),
		(x"38fe197ebf9407fa00f2a6ec8d47fa00", x"1e4dc5d24b75b8a1", x"254CAB64F613CA71"),
		(x"733ccd6f3f79c1d853601f0c53346d6a", x"5df367829ff0e2f3", x"0D0EDFB2D807B32C"),
		(x"8acc2aa266cbbe843b51f8d6fb14612a", x"a957a0fed8d56b5e", x"C4E2E776935198D4"),
		(x"b310922cc6f2e41d004ac89349f37d62", x"ef86492cce0469a6", x"BCE881F6EC785F86"),
		(x"baf9621f6b5f79dcac1a65c73e44740d", x"ca7292cbec11f9fa", x"EE9BBDE6F36844BE"),
		(x"9209a3f916c68f187d1f0295af33d816", x"7f39cc7b52775bba", x"D0BD7A90C725E785"),
		(x"7f77ea3931afe959cd52a9e0c85a1b23", x"b010d57459116b01", x"3126AEC88413CD2F"),
		(x"d0498a7581b2f15d5ffc9e894648e493", x"277c121f122ef5fa", x"821FF4930F95F8FD"),
		(x"2040f1f7279ebcaa3b9583e77a6ebb60", x"2bc24c9d44548236", x"D71C9C0DEC2D1A76"),
		(x"783e5138eb33ec8b56c025ad3482bfb9", x"9f57caf7a60d3e02", x"0B55EEF26D20C797"),
		(x"f3d6d17252bc3dca89d3067844a64b4b", x"ce32f7ca58a2a4a8", x"12C5419C5BAB2633"),
		(x"ba6b9780a172f6f7ecadb1f3500bddb7", x"bd9f4d7c9f85b718", x"855B0CEDB81DF9EE"),
		(x"2ab751328f99c7653e4c1de267cac34d", x"6aeca5a1dafc1c3e", x"85BD3FF44018F631"),
		(x"97282802bdee742b93996eab855b8bd5", x"c8f3cfce121d5e88", x"FB69E92B57588AFF"),
		(x"c3c0735abd74d4826cf6a524d588bc60", x"8142f5650893f6e7", x"97E9FBC28F90DDF3"),
		(x"68c49f9139eff7190ad61e717ff19ece", x"ef2934bab53bd298", x"2419CBDF392DC108"),
		(x"ab6490d306c0f2cf150a4270b3f6fd27", x"93f9f6588c5e634a", x"F07DE481014AEFD2"),
		(x"a7f049c2e4f1618362bfa60e3dcc5909", x"827449b14041b156", x"9F0B585FE66BFE63"),
		(x"56647b7ce995d93605509d6ee919445e", x"5d414d71f4f15fb8", x"7872AE571BDB6E2A"),
		(x"59dc4270e3630f5cffc1f1708f5efb34", x"f8591a104fbb4293", x"645DDC4CBDC60A29"),
		(x"274ad3af59087f8d5d3877d7e8fdf778", x"6ae8b76bc8ddcfd0", x"DF6805FD50F31C23"),
		(x"cc618f69f481e33f6940d030c0be35eb", x"9503c32438e7b9a2", x"538CF04F4B46A4BC"),
		(x"645279e1ac1a07adc47e5f2e452d2771", x"59018eb8ab49f069", x"42B48A8056B06A76"),
		(x"39c37eed4d0610adb51fc9d6beb7c026", x"e5582e08ff58e0bc", x"E7992D832AB0834D"),
		(x"743f2b0d60085f7e7ab4092b8a707706", x"c06b1dd465b065f7", x"0FAE480CE2A657B6"),
		(x"e268779ef74b1addf3ce84567a7c3c41", x"5560ed5aeb6970d7", x"5B9F561AD8D9028E"),
		(x"e2cb1a91d4b3874eec675a90bc701e36", x"752e3b89a5e114e0", x"2AC16EBD2224A9C9"),
		(x"707b0ddd8c8d251c2142ec05712fa835", x"8dae77cd7a2b4659", x"4ED98BF51939C225"),
		(x"98c668a7d4aff4f170cf4e600315740c", x"1538290581dcb984", x"7F7EEF63DE351181"),
		(x"98bce3cc892322be53c66af92f9c910a", x"22b9e246fbd95439", x"7A0508A9140B4428"),
		(x"d383dccd44cfcb1d5cb4c9f5afd898d9", x"3b9987f0336a9e59", x"A649243F852C66B6"),
		(x"36365c593b7df2c053ccb74d71c562f6", x"acb30a09a8178961", x"3AC7DA9BAA913EF3"),
		(x"09820404d77964cd200ce894f070fd6d", x"1adc9d4f125ed5b5", x"06103ECD7A0938C3"),
		(x"1d8e4d33dfc1232ed9030409801404ea", x"ef426eb4484a6ccf", x"201C43CC60B51D23"),
		(x"481de2bec525007c53ea855dcbf7e484", x"90a54b32f4c3a956", x"CD18AF79DFAE24D6"),
		(x"ecd1bec787bb11e92e1a2d041c7a481f", x"15b6e5d46d71cc5d", x"7BFA6E1A43E951E9"),
		(x"0ef6beb19f28aa12c61bfa63117510f4", x"4a2ffd8f14424c6f", x"009B67D47A16C59A"),
		(x"c40ca33cb8e36ae973cd2b414d845531", x"7976930299b787d2", x"68AA18778001CCD9"),
		(x"855dd59bc428a065bc8d8429294d450a", x"00e1bd6eeb86747c", x"EBDE32E33CEC7D07"),
		(x"34f1c14b3ebec303e0f117c3a8acd818", x"6a7bbd1510dc9053", x"E66A30605929B36D"),
		(x"756f3fc0a5b58d8d5cabaec132c0f065", x"5606daf6b9c19184", x"109949E883FFEF14"),
		(x"6d2d1d27b044810284d8de60d94df1d2", x"bd3ce81327872fde", x"796E22F38F52B160"),
		(x"bb01e74f4ea6b9a8b2609422fedd4c4a", x"0a01b3ea9d20a822", x"CCA1096B05E0FF80"),
		(x"ed1300cc430f413262190dea4607ac0c", x"01309043b31036fc", x"0BD189666F5650AE"),
		(x"a8cfb2cfabac0ef91f837d584857ce90", x"63e05b8673ed2c6c", x"E286F319BCE79937"),
		(x"caeaadc532fa605c7595d800a468f47b", x"70f814e97367733a", x"064A01E41829B167"),
		(x"9addf440bda1ff69fab0e97db30d77f5", x"36853b86d9526904", x"FBFE06A4624C2F9E"),
		(x"bfa40918e511c53a5923301de0db4d96", x"0f89d28ac337c751", x"9F9EA16EECF20797"),
		(x"10d94467d7df52adfb787bbb3b03c45b", x"ba223e0d44c297d7", x"BF48AF540875BADA"),
		(x"ebfa8e9b19f70a7ffc8ce84ae9b42149", x"d7b3caec00a1fbe1", x"0DB30A4533E8E266"),
		(x"65cd1f847413aa835d0a549bd629d046", x"28faaa04735925c1", x"7049BD1521D28D26"),
		(x"2f01e822541953f8264cda876c1cabc8", x"7d360b1c0592e8ed", x"91B6851AF086E5BA"),
		(x"703c08217aa8e10119027fc249ec5ddc", x"00f8b3bec170bdea", x"77DEC679EB14B509"),
		(x"bd046beb19b6fb531ff12b089294c7b6", x"074bf36e00742947", x"06C544A56719EBB3"),
		(x"c697e5703cb170bd4d11c77c3659fa73", x"a0f96ade8e9bf2e0", x"C638B82FBD7913B2"),
		(x"0423a7000553df2f508c0fb3eeadf3c5", x"cce9e546ce7aa82c", x"A67B4B31304BCAF9"),
		(x"df0a959a770370e032e30d65d18babd5", x"c8e2af95f14c23c8", x"E411936126E39A98"),
		(x"ec09bd9ccb663b12fff4fbb1e926bb56", x"2f26409bee5bc3e9", x"7F33107BFF75C65B"),
		(x"01f0d72c88043b3779b476e69966afbd", x"5f3d0f7158767ea8", x"0F3D2953649DF139"),
		(x"c65a9ffe42988c6ac851f1996dea7e6c", x"dc1b35440693437b", x"3AE2B263B7CBE303"),
		(x"8b3bfd57b831da2bde9b4625750c59e5", x"cfe04377b599c5da", x"43B2B932320C28CF"),
		(x"72d02559d3641c4436e2792336f26bea", x"51fc54604145a48a", x"5A7F7656262B225E"),
		(x"4a916c73b14da0a61e262344220e0140", x"911195998be342fa", x"AC17D57D665A711F"),
		(x"27521f6714ab7d28a058c8b91f385483", x"9b66843f786d851a", x"AD87DA0740F80408"),
		(x"20c9d53e8c377e1d79b954c895c89358", x"16c921e5e9ee84b8", x"8DE9C56D7CF9E283"),
		(x"781954a7fbd52ea1b84267b1169aeee4", x"48f7d37a36001eb3", x"0558EF640823F788"),
		(x"a3ec65cdd6632747a45f913d3b1b3a8b", x"31485a12e1e3a9c3", x"3F64B0A4724144AE"),
		(x"7ec1175e47d862deba22e94f4206b40b", x"1fceba4edccd2b46", x"4A49BC2F8EB55790"),
		(x"463ac1751ee568cebf858299388f0060", x"6fc214208d319ad3", x"815D3DB1E6183E65"),
		(x"9aed37f37783c2d0ea77472ce7358cf4", x"b89db8a5e0d0a207", x"4069F625149C072C"),
		(x"7f55a833153f80e3fb19117bba8e99ae", x"a8c8ff69d872b574", x"F9C307A88F907F7C"),
		(x"37404b7a6ef1d0b2e4d573d5385591bc", x"0aa57bed7a504f81", x"FEF1994D8FC65257"),
		(x"662cbdde6d5ad23bcd16d0e723a2f76d", x"f6883e025dcce06d", x"3E33E89B8141B009"),
		(x"76f214b926b6990293123b8013c84d9b", x"d937843eec3a56bb", x"D6CEAE83DE53521B"),
		(x"c7cb186148797db6963e903b74db2c0a", x"22ae9195d0047c6e", x"1B808FDDA6B8932A"),
		(x"03a7a290bdf7c2627a1f7a6240fd36d7", x"08bfe5e3c1308af2", x"B597F2B7B27BB58C"),
		(x"0eecb149ff7b74cda548ec855fe1f534", x"9d4bbafb624ad73a", x"35C72C7803ED793A"),
		(x"e6a8184146e92ff6ddb6955ce9485939", x"af5a1dbe7c62b7ae", x"EF6FA30DFD80AB28"),
		(x"e7db178d3f4d519ec3ce6509f5316958", x"b272a3b85251ad00", x"27CB522596146E46"),
		(x"2d940db5c7ea54a521499afa8ad57354", x"71e39c3fa60c38bd", x"940D822AD08AF191"),
		(x"e72d83b3b280b03371b59c3f78ce4367", x"32455ae9a4cfcd2a", x"6DE2D9E31C956665"),
		(x"61a490af1e6fc8332761d7123cb1fdeb", x"89e0cad555e15e4b", x"92299C7B24EBB067"),
		(x"ff632111151af03cdd28baa40cbdf387", x"6232b0c367cb4d7e", x"EE1D61220C07D9F8"),
		(x"670e1de29a5c810edf2dfdc01f2f2b6f", x"7e551b30fa6d1dd1", x"8CC2292F360CEF79"),
		(x"71537f5fee2a8ad81592af014833d1c0", x"bb31a4956373bd23", x"4B6EE33767C0D231"),
		(x"25c4b9cdfa0f1e9e7997b3d9b06fad98", x"25aefb1a625ec374", x"180C5A2F0E228B9E"),
		(x"954e3b31979fc83c1a63e0b011e8cc08", x"b2f188112082e050", x"D30A21E71F544DE2"),
		(x"e63b20f08f5a757bf25e6fa500e5fcdd", x"0611c0a6446e1006", x"CF3D94E44CD4F13D"),
		(x"7bfda3d7016723518fde184667c424ff", x"c54fb189cce1f91a", x"9096643ECF86EB26"),
		(x"8388e211040eaecbef10ca0331462bac", x"c3227b69ed81b62e", x"3A00071BDE5D2066"),
		(x"288cafbfd571e8244cd67ff21d01ca1f", x"1322ddf4752c1f8d", x"62531DC2FE930F44"),
		(x"2c4c763709e16ee8ba4f5e77e141cf69", x"8b4e02ec304a3f9e", x"87385BC86FEBE649"),
		(x"26bb07a04fff921428892ef486e09738", x"4bf7b7e5296d89a4", x"6C8390025A563EA8"),
		(x"959e4a300b219c65652094297ab7a690", x"be60310ddafd218b", x"8EBB9A1926F15F41"),
		(x"1fdece37ab5653c5e0170fcf21dbab43", x"f8efafb7136688a7", x"D162824F825936D6"),
		(x"f592fb6c157554a3ec5e27b62b6c707b", x"6055fac8b9a88dea", x"F8105A7F8FBBB56C"),
		(x"6f1fd2ef2a11f5fe4075203aee79c1d0", x"1ec456dbc8d6a214", x"A481F8B80367E0B7"),
		(x"f8445282e9c86dbbfbf3982f7f774343", x"4c1f2d9fcc76d8ff", x"F54C618DABC0E7F9"),
		(x"c2cffd00fa2b6919c2da298d7a83c4ab", x"8249f236cb2a697a", x"E460B1B9FABA0740"),
		(x"21b45543f49151a98d225abf4358ad21", x"0ea217ca8fcf6620", x"FA657E4C862930B3"),
		(x"b7bb96bec7a27725989c45935ea7cf9c", x"ae8182ef4f5d77d8", x"A9391DAB5382AA4A"),
		(x"855cd27039d321a773d155c508cec6a3", x"76b1ba1504b7e5e7", x"329A06F00EAD8B87"),
		(x"2c43fb6997d68dccb2833261ac0d7a7b", x"1ef1e2384704ade1", x"3910E528788E3161"),
		(x"760fdd83795f72bfc5ea82700aa26f7e", x"fd997dda51321d26", x"9EC5B3C22752F4F5"),
		(x"07e136fd04dab231ad31ceb1dad08f25", x"30df6960ebaf5a5b", x"5F7471ECB475DD9D"),
		(x"56fe73cdc65f8f03ee549dc8f4e47e8b", x"cb5c8eeee8e2b530", x"95939C91931B0473"),
		(x"ac7619cc99d9bcfbffe80197f37f9221", x"4cfe6da0df40307f", x"4B91EF59425CA2BB"),
		(x"0831a47a84061240d6de2ba647efdd0e", x"ec4ed4eea382a9e5", x"AC8E6FF4A94CD0AC"),
		(x"45654063e150cbb0a97ce6d48fb9e727", x"d7681c2d27585daf", x"D3750B279FE26267"),
		(x"4605f9e37883e0b3d8eadff0c67f0cd5", x"88177cd1f644e714", x"C0C557B125FE3BBB"),
		(x"a33233a5f2c2f06b3f51b09ea8f21d8e", x"3f9f74a7b9c0e1b2", x"DC519A6356C3BB74"),
		(x"6d117d4a2b8cdc58b6a5d1a850de3a0e", x"e0655ea10a0f4578", x"9D2683DBC2468B1C"),
		(x"b6a6ee8109ae015b81804d3cc713268e", x"7fe9da24ac8aa1b2", x"9BA60D7D23DAE715"),
		(x"ad6fd0b86775cbe2e3d4432696f65944", x"d428084ca75cf4b8", x"ED51D1640D9B71E4"),
		(x"568982c94a430fd975e5aa0b52d5e43b", x"e7a79a33e14abc8e", x"0C4AFC52CD17EB88"),
		(x"17c7e47e73ca3167335c58e4d5dc4799", x"487297324fd1e332", x"0B5C5AB4E156DA21"),
		(x"12f500f105d3b1a8499ea920b40941ce", x"d75edc50fba3f005", x"62CD1D6FA67278F7"),
		(x"29a637f8e671dd74dcd92c2e2ae394cc", x"d3dc6146e92b3b10", x"35E3A25228EB74EB"),
		(x"575bd4bfdf8c8022761908dfcf029a59", x"44bb6b2340576a49", x"C168E9350C8684B9"),
		(x"4d9bc7f20e36e530dcb1b4567fb46b80", x"a48568ae9ef3abe2", x"B4ED571659DCE957"),
		(x"62ad435a0ce0083cb71e84ec09eff7c0", x"dd8f5c7a80cc7af1", x"55D9A84B9F07C836"),
		(x"81c4f6deffb07647f8cabea916a035ad", x"bb5fc7f0dd315be1", x"7645398005F706DA"),
		(x"e5e02b030ec3e7ad7088b71e70844b82", x"9ee57c53988192de", x"E2A2D8891C9E94CE"),
		(x"adbd8726f65bcc9fec7bcabafe6d5a00", x"5de43c3177dd5b52", x"62971F070E79775F"),
		(x"4bef944323249841f4cdb3d97f9a6ae3", x"9eb5cb3ff811fd58", x"7F1750C69547D8BE"),
		(x"065170186580bca6b42b0103bf3490c1", x"d209739a1a0d3f72", x"DFA92B6B6E13DC36"),
		(x"136e25a6175da08e609dfbd62ee26a94", x"acc2ac2b1ca235a0", x"3CBE87236CFC57B1"),
		(x"8e9be09c46b91f8602b8aa9c611408da", x"5a869fda9262905b", x"D83BCC56291EF05C"),
		(x"9affa7384f026af9174d8025d11bc780", x"da9535abd54a149e", x"E4D601504A4D741E"),
		(x"4af7b74c30ae71d829428dc594964390", x"0a83143737028ffa", x"ABDF6A90FA5B5E2D"),
		(x"2c22e009a14239baacf2fcfc0ff3ee20", x"a13c2ad485c69f5e", x"681F7B215E96217E"),
		(x"5525126e8af6b513131350797f805b9d", x"cc0a69c315f2d18f", x"0ADA061CB652F43B"),
		(x"b3f3cf367a2a9c16396e4d562a3768de", x"82ca9cc3f222da7c", x"796FEB91AEB0F0AF"),
		(x"0d1271bb0e7858a2db882b50963561b9", x"e57eeeef26de39be", x"9A9E42CF6871FA38"),
		(x"3d0f6639f8b6127ab5ca89845417a19c", x"43891b72c85cfb86", x"2CC37BB585357D47"),
		(x"fc06891eb1712620efab5340bea84555", x"2555733d13bf8f05", x"EBE7FEF5A5D2E4E7"),
		(x"5691ccc74db94d095b47f043e703003f", x"aa6b79ebcf9c7533", x"D6EC73982012CE5C"),
		(x"b9f945a718e9b9a6fe427f8a420d2c33", x"4084c1022148d45a", x"BABF044F2E0505FF")
    	);
end package prince_cipher_pkg;


